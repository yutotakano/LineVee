module linevee
